Hi & Welcome to the Program , 
 This program is a collection of the capabilities of using the Registery 
To Get Data about Your PC and Writing Data Again, 
It Conatins The Following : 
1) Special Folder's Path's : ( ONLY  5 LINES OF CODE )
( 'Desktop' , 'Programs' , 'Favorites' , 'History' ,Administrative Tools;   AppData;cookies;desktop;favorites
;fonts;history;Local AppData;Local settings;my music;my pictures
 my vedio;nethood;personal;printhood;programs;recent;send to;start menu;startup;templates)
		
 2)The Previous Keywords Used in Search , This words can't be removed , 
     Now You can Remove it Very Easy or even replace it , 

3) The History of URL Visited , You can remove only one or two URLs or whatever  without Loosing the Rest , 

4) Changing the HomePage ,
 
ALL THAT WITHOUT ANY API'S  , A  FREE  API  CODE .

****** NO One LINE OF API IS USED*************